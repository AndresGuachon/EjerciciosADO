----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    08:22:37 05/24/2022 
-- Design Name: 
-- Module Name:    Ej1_17 - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity Ej1_17 is
    Port ( a0, b0 : in  STD_LOGIC;
           a1, b1 : in  STD_LOGIC;
           a2, b2 : in  STD_LOGIC;
           a3, b3 : in  STD_LOGIC;
           F : out  STD_LOGIC);
end Ej1_17;

architecture Behavioral of Ej1_17 is

begin


end Behavioral;

