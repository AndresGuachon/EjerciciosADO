----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    08:31:15 05/24/2022 
-- Design Name: 
-- Module Name:    Ej1_21 - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity Ej1_21 is
    Port ( botonA, botonB : in  STD_LOGIC;
           giro : out  STD_LOGIC);
end Ej1_21;

architecture Behavioral of Ej1_21 is

begin
		process(botonA, botonB)
		begin
			if(botonA='1') then giro <='1';
			elsif (botonB = '1') then giro <='0';
			end if;
			end process;


end Behavioral;

