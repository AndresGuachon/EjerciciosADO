----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    08:18:30 05/24/2022 
-- Design Name: 
-- Module Name:    Ej1_11_2 - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity Ej1_11_2 is
    Port ( A : in  STD_LOGIC_VECTOR (0 downto 3);
           B : in  STD_LOGIC_VECTOR (0 downto 3);
           C : out  STD_LOGIC_VECTOR (0 downto 3));
end Ej1_11_2;

architecture Behavioral of Ej1_11_2 is

begin


end Behavioral;

